`include "define.v"
module ex(
    input wire rst,
    //译码阶段传递过来的操作码及数据
    input wire [`AluOpBus]      aluop_i,
    input wire [`AluSelBus]     alusel_i,
    input wire [`RegBus]        reg1_i,
    input wire [`RegBus]        reg2_i,
    input wire [`RegAddrBus]    wd_i,
    input wire                  wreg_i,

    //执行的结果
    output reg[`RegAddrBus]     wd_o,
    output reg[`RegBus]         wdata_o,
    output reg                  wreg_o,

	//从hilo_reg模块传递过来的数据
	input wire [`RegBus] 		hi_i,
	input wire [`RegBus] 		lo_i,
	//位于访存阶段对hilo_reg寄存器读写情况
	input wire 					mem_whilo_i,
	input wire [`RegBus] 		mem_hi_i,
	input wire [`RegBus] 		mem_lo_i,
	//位于回写阶段对hilo_reg寄存器的读写情况
	input wire	 				wb_whilo_i,
	input wire [`RegBus] 		wb_hi_i,
	input wire [`RegBus] 		wb_lo_i,
	
	//对寄存器修改情况的输出
	output reg					whilo_o,
	output reg [`RegBus] 		hi_o,
	output reg [`RegBus] 		lo_o,
	
	//多周期执行性指令控制
	input wire [`DoubleRegBus]	hilo_temp_i,
	input wire [1:0] 			cnt_i,
	output reg [`DoubleRegBus]  hilo_temp_o,
	output reg [1:0] 			cnt_o,
	output reg 					stallreq_from_ex,
	
	//除法指令新增信号
	input wire [`DoubleRegBus] 	div_result_i,
	input wire 					div_ready_i,
	output reg 					signed_div_o,
	output reg [`RegBus] 		div_opdata1_o,
	output reg [`RegBus] 		div_opdata2_o,
	output reg 					div_start_o,
	
	//转移指令
	input wire 					is_in_delayslot_i,
	input wire [`RegBus] 		link_address_i,
	
	//加载存储指令
	input wire [`RegBus] 		inst_i,
	output wire [`AluOpBus] 	aluop_o,
	output wire [`RegBus] 		mem_addr_o,
	output wire [`RegBus]       reg2_o
	
);

assign aluop_o=aluop_i;
assign mem_addr_o=reg1_i+{{16{inst_i[15]}},inst_i[15:0]};
assign reg2_o=reg2_i;

reg [`RegBus]   logicount;		//
reg [`RegBus]  	shiftres;		//
reg [`RegBus]   moveres;		//
reg [`RegBus]  	HI; 			//
reg [`RegBus]  	LO;				//
reg [`DoubleRegBus] 	mulres;	//
reg [`RegBus]  	arithmeticres;	//

wire 			ov_sum;			//
wire [`RegBus] 	result_sum;		//
wire [`RegBus] 	reg2_i_mux;		//
wire 			reg1_lt_reg2;	//
wire [`RegBus] 	reg1_i_not;  	//

wire [`RegBus] opdata1_mux;  	//
wire [`RegBus] opdata2_mux;  	//
wire [`DoubleRegBus] hilo_temp;	   //
reg  [`DoubleRegBus] hilo_temp1;
reg  				 stallreq_for_madd_msub;

reg 			stallreq_for_div;


//有符号加法运算或减法运算数据处理
assign reg2_i_mux=((aluop_i==`EXE_SUB_OP)||(aluop_i==`EXE_SUBU_OP)
					||(aluop_i==`EXE_SLT_OP))?(~reg2_i+1'b1):reg2_i; 
assign result_sum=reg1_i+reg2_i_mux;
assign ov_sum=((!reg1_i[31])&&(!reg2_i_mux[31])&&result_sum[31])
				||(reg1_i[31]&&reg2_i_mux[31]&&(!result_sum[31]));
//判断reg1<reg2
assign reg1_lt_reg2=(aluop_i==`EXE_SLT_OP)?((reg1_i[31]&&(!reg2_i[31]))||(!reg1_i[31]&&!reg2_i[31]&&result_sum[31])
											||(reg1_i[31]&&reg2_i[31]&&result_sum[31])):(reg1_i<reg2_i);
assign reg1_i_not=~reg1_i;

//有符号乘法运算数据处理
assign opdata1_mux=(((aluop_i==`EXE_MUL_OP)||(aluop_i==`EXE_MULT_OP)||(aluop_i==`EXE_MADD_OP)||(aluop_i==`EXE_MSUB_OP))&&reg1_i[31])?(~reg1_i+1'b1):reg1_i;
assign opdata2_mux=(((aluop_i==`EXE_MUL_OP)||(aluop_i==`EXE_MULT_OP)||(aluop_i==`EXE_MADD_OP)||(aluop_i==`EXE_MSUB_OP))&&reg2_i[31])?(~reg2_i+1'b1):reg2_i;
assign hilo_temp=opdata1_mux*opdata2_mux;

//简单算术运算				
always @(*) begin
	if(rst==`RstEnable) begin
		arithmeticres<=`ZeroWord;
	end else begin
		case(aluop_i)
			`EXE_ADD_OP,`EXE_ADDU_OP,`EXE_ADDI_OP,`EXE_ADDIU_OP: begin
				arithmeticres<=result_sum;
			end
			`EXE_SLT_OP,`EXE_SLTU_OP: begin
				arithmeticres<=reg1_lt_reg2;
			end
			`EXE_SUB_OP,`EXE_SUBU_OP: begin
				arithmeticres<=result_sum;
			end
			`EXE_CLZ_OP: begin
				arithmeticres<=reg1_i[31]?0:reg1_i[30]?1:reg1_i[29]?2
							   :reg1_i[28]?3:reg1_i[27]?4:reg1_i[26]?5
							   :reg1_i[25]?6:reg1_i[24]?7:reg1_i[23]?8
							   :reg1_i[22]?9:reg1_i[21]?10:reg1_i[20]?11
							   :reg1_i[19]?12:reg1_i[18]?13:reg1_i[17]?14
							   :reg1_i[16]?15:reg1_i[15]?16:reg1_i[14]?17
							   :reg1_i[13]?18:reg1_i[12]?19:reg1_i[11]?20
							   :reg1_i[10]?21:reg1_i[9]?22:reg1_i[8]?23
							   :reg1_i[7]?24:reg1_i[6]?25:reg1_i[5]?26
							   :reg1_i[4]?27:reg1_i[3]?28:reg1_i[2]?29
							   :reg1_i[1]?30:reg1_i[0]?31:32;
			end
			`EXE_CLO_OP: begin
				arithmeticres<=reg1_i_not[31]?0:reg1_i_not[30]?1:reg1_i_not[29]?2
							   :reg1_i_not[28]?3:reg1_i_not[27]?4:reg1_i_not[26]?5
							   :reg1_i_not[25]?6:reg1_i_not[24]?7:reg1_i_not[23]?8
							   :reg1_i_not[22]?9:reg1_i_not[21]?10:reg1_i_not[20]?11
							   :reg1_i_not[19]?12:reg1_i_not[18]?13:reg1_i_not[17]?14
							   :reg1_i_not[16]?15:reg1_i_not[15]?16:reg1_i_not[14]?17
							   :reg1_i_not[13]?18:reg1_i_not[12]?19:reg1_i_not[11]?20
							   :reg1_i_not[10]?21:reg1_i_not[9]?22:reg1_i_not[8]?23
							   :reg1_i_not[7]?24:reg1_i_not[6]?25:reg1_i_not[5]?26
							   :reg1_i_not[4]?27:reg1_i_not[3]?28:reg1_i_not[2]?29
							   :reg1_i_not[1]?30:reg1_i_not[0]?31:32;
			end
			default: begin
			end
		endcase			
	end
end
//乘法运算结果
always @(*) begin
	if(rst==`RstEnable) begin
		mulres<={`ZeroWord,`ZeroWord};
	end else if((aluop_i==`EXE_MULT_OP)||(aluop_i==`EXE_MUL_OP)
				  ||(aluop_i==`EXE_MADD_OP)||(aluop_i==`EXE_MSUB_OP)) begin
		if(reg1_i[31]^reg2_i[31]==1'b1) begin
			mulres<=~hilo_temp+1'b1;
		end else begin
			mulres<=hilo_temp;
		end
	end else begin
		mulres<=hilo_temp;
	end
end

//madd,maddu,msub,msubu指令
always @(*) begin
	if(rst==`RstEnable) begin
		hilo_temp_o<={`ZeroWord,`ZeroWord};
		cnt_o<=2'b00;
		stallreq_for_madd_msub<=`NoStop;
	end else begin
		case(aluop_i)
			`EXE_MADD_OP,`EXE_MADDU_OP: begin
				if(cnt_i==2'b00) begin
					hilo_temp_o<=mulres;
					cnt_o<=2'b01;
					hilo_temp1<={`ZeroWord,`ZeroWord};
					stallreq_for_madd_msub<=`Stop;
				end else if(cnt_i==2'b01) begin
					hilo_temp_o<={`ZeroWord,`ZeroWord};
					cnt_o<=2'b10;
					hilo_temp1<=hilo_temp_i+{HI,LO};
					stallreq_for_madd_msub<=`NoStop;
				end
			end
			`EXE_MSUB_OP,`EXE_MSUBU_OP: begin
				if(cnt_i==2'b00) begin
					hilo_temp_o<=~mulres+1'b1;
					cnt_o<=2'b01;
					hilo_temp1<={`ZeroWord,`ZeroWord};
					stallreq_for_madd_msub<=`Stop;
				end else if(cnt_i==2'b01) begin
					hilo_temp_o<={`ZeroWord,`ZeroWord};
					cnt_o<=2'b10;
					hilo_temp1<=hilo_temp_i+{HI,LO};
					stallreq_for_madd_msub<=`NoStop;
				end
			end
			default: begin
				hilo_temp_o<={`ZeroWord,`ZeroWord};
				cnt_o<=2'b00;
				stallreq_for_madd_msub<=`NoStop;
			end
		endcase
	end
end
always @(*) begin
	stallreq_from_ex=stallreq_for_madd_msub||stallreq_for_div;
end

//除法运算
always @(*) begin
	if(rst==`RstEnable) begin
		stallreq_for_div<=`NoStop;
		div_opdata1_o<=`ZeroWord;
		div_opdata2_o<=`ZeroWord;
		div_start_o<=`DivStop;
		signed_div_o<=1'b0;
	end else begin
		stallreq_for_div<=`NoStop;
		div_opdata1_o<=`ZeroWord;
		div_opdata2_o<=`ZeroWord;
		div_start_o<=`DivStop;
		signed_div_o<=1'b0;
		case(aluop_i) 
			`EXE_DIV_OP:	begin
				if(div_ready_i==`DivResultNotReady) begin
					stallreq_for_div<=`Stop;
					div_opdata1_o<=reg1_i;
					div_opdata2_o<=reg2_i;
					div_start_o<=`DivStart;
					signed_div_o<=1'b1;
				end else if(div_ready_i==`DivResultReady) begin
					stallreq_for_div<=`NoStop;
					div_opdata1_o<=reg1_i;
					div_opdata2_o<=reg2_i;
					div_start_o<=`DivStop;
					signed_div_o<=1'b1;
				end else begin
					stallreq_for_div<=`NoStop;
					div_opdata1_o<=`ZeroWord;
					div_opdata2_o<=`ZeroWord;
					div_start_o<=`DivStop;
					signed_div_o<=1'b0;
				end
			end
			`EXE_DIVU_OP:	begin
				if(div_ready_i==`DivResultNotReady) begin
					stallreq_for_div<=`Stop;
					div_opdata1_o<=reg1_i;
					div_opdata2_o<=reg2_i;
					div_start_o<=`DivStart;
					signed_div_o<=1'b0;
				end else if(div_ready_i==`DivResultReady) begin
					stallreq_for_div<=`NoStop;
					div_opdata1_o<=reg1_i;
					div_opdata2_o<=reg2_i;
					div_start_o<=`DivStop;
					signed_div_o<=1'b0;
				end else begin
					stallreq_for_div<=`NoStop;
					div_opdata1_o<=`ZeroWord;
					div_opdata2_o<=`ZeroWord;
					div_start_o<=`DivStop;
					signed_div_o<=1'b0;
				end
			end
			default:	begin
			end
		endcase
	end
end


//读取HI和LO寄存器内的值
always @(*) begin
	if(rst==`RstEnable) begin
		HI<=`ZeroWord;
		LO<=`ZeroWord;
	end else if(mem_whilo_i==`WriteEnable) begin
		{HI,LO}<={mem_hi_i,mem_lo_i};
	end else if(wb_whilo_i==`WriteEnable) begin
		{HI,LO}<={wb_hi_i,wb_lo_i};
	end else begin
		{HI,LO}<={hi_i,lo_i};
	end
end
//移动操作指令执行
always @(*) begin
	if(rst==`RstEnable) begin
		moveres<=`ZeroWord;
	end else begin
		moveres<=`ZeroWord;
		case(aluop_i)
			`EXE_MFHI_OP: 	begin
				moveres<=HI;
			end
			`EXE_MFLO_OP: 	begin
				moveres<=LO;
			end
			`EXE_MOVN_OP: 	begin
				moveres<=reg1_i;
			end
			`EXE_MOVZ_OP:	begin
				moveres<=reg1_i;
			end
			default:	begin
			end
		endcase
	end
end
//写HI和LO寄存器操作
always @(*) begin
	if(rst==`RstEnable) begin
		whilo_o<=`WriteDisable;
		hi_o<=`ZeroWord;
		lo_o<=`ZeroWord;
	end else if((aluop_i==`EXE_DIV_OP)||(aluop_i==`EXE_DIVU_OP)) begin
		whilo_o<=`WriteEnable;
		hi_o<=div_result_i[63:32];
		lo_o<=div_result_i[31:0];
	end else if((aluop_i==`EXE_MSUB_OP)||(aluop_i==`EXE_MSUBU_OP)) begin
		whilo_o<=`WriteEnable;
		hi_o<=hilo_temp1[63:32];
		lo_o<=hilo_temp1[31:0];
	end else if((aluop_i==`EXE_MADD_OP)||(aluop_i==`EXE_MADDU_OP)) begin
		whilo_o<=`WriteEnable;
		hi_o<=hilo_temp1[63:32];
		lo_o<=hilo_temp1[31:0];
	end else if((aluop_i==`EXE_MULT_OP)||(aluop_i==`EXE_MULTU_OP)) begin
		whilo_o<=`WriteEnable;
		hi_o<=mulres[63:32];
		lo_o<=mulres[31:0];
	end else if(aluop_i==`EXE_MTHI_OP) begin
		whilo_o<=`WriteEnable;
		hi_o<=reg1_i;
		lo_o<=LO;
	end else if(aluop_i==`EXE_MTLO_OP) begin
		whilo_o<=`WriteEnable;
		hi_o<=HI;
		lo_o<=reg1_i;
	end else begin
		whilo_o<=`WriteDisable;
		hi_o<=`ZeroWord;
		lo_o<=`ZeroWord;
	end	
end


//依据aluop_i的数据进行指令操作，逻辑运算指令
always @(*) begin
    if(rst==`RstEnable) begin
        logicount<=`ZeroWord;
    end else begin
        case(aluop_i)
            `EXE_OR_OP: begin
                logicount<=reg1_i|reg2_i;
            end
			`EXE_AND_OP: begin
				logicount<=reg1_i&reg2_i;
			end
			`EXE_NOR_OP: begin
				logicount<=~(reg1_i|reg2_i);
			end
			`EXE_XOR_OP: begin
				logicount<=reg1_i^reg2_i;
			end
            default: begin
                logicount<=`ZeroWord;
            end
        endcase
    end
end

//根据aluop_i进行指令操作，移位运算符
always @(*) begin
	if(rst==`RstEnable) begin
		shiftres<=`ZeroWord;
	end else begin
		case(aluop_i)
			`EXE_SLL_OP: begin
				shiftres<=reg2_i<<reg1_i[4:0];
			end
			`EXE_SRL_OP: begin
				shiftres<=reg2_i>>reg1_i[4:0];
			end
			`EXE_SRA_OP: begin
				shiftres <=({32{reg2_i[31]}}<<(6'd32-{1'b0,reg1_i[4:0]}))|reg2_i>>reg1_i[4:0];
			end
			default: begin		
				shiftres<=`ZeroWord;
			end
		endcase
	end
end


//根据alusel_i指示的运算类型选择最终运算结果
always @(*) begin
    wd_o<=wd_i;
	if(((aluop_i==`EXE_ADD_OP)||(aluop_i==`EXE_ADDI_OP)||(aluop_i==`EXE_SUB_OP))&&(ov_sum==1'b1)) begin
		wreg_o<=`WriteDisable;
	end else begin
		wreg_o<=wreg_i;
	end
    case(alusel_i)
        `EXE_RES_LOGIC: begin
            wdata_o<=logicount;
        end
		`EXE_RES_SHIFT: begin
			wdata_o<=shiftres;
		end
		`EXE_RES_MOVE: 	begin
			wdata_o<=moveres;
		end
		`EXE_RES_ARITHMETIC: begin
			wdata_o<=arithmeticres;
		end
		`EXE_RES_MUL: begin
			wdata_o<=mulres[31:0];
		end
		`EXE_RES_JUMP_BRANCH:	begin
			wdata_o<=link_address_i;
		end
        default: begin
            wdata_o<=`ZeroWord;
        end
    endcase
end

endmodule 
